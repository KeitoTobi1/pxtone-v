module pxtone

struct Pxtone {
	core C.MPXTN
}

pub fn pxtone_load(){

}

pub fn pxtone_start(){

}