module pxtone

struct Pxtone {
	core Mpxtn
}

pub fn pxtone_load(){

}

pub fn pxtone_start(){

}