module pxtone

struct Pxtone {}

pub fn pxtone_load(){

}

pub fn pxtone_start(){

}