module pxtone

const (
	EVENT_MAX = 50000
	MPXTN_SPS = 44100
	MPXTN_BPS = 8
	MPXTN_CH = 2
	FILESIZE_MAX = (32*1024*1024)
	VOL_MAX = 128
	PAN_MAX = 128
)